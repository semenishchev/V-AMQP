module main
// import vamqp

fn main() {
	println('Hello World!')
}
