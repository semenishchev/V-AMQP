module vamqp

struct Delivery { // TODO: fill the struct

}