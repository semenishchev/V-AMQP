module vamqp

fn main() {
	println('Hello World!')
}
